module counter #(
    parameter WIDTH = 8
)(
    // Interface signals
    input logic clk,                // clock
    input logic rst,                // reset
    input logic en,                 // load counter from data
    output logic [WIDTH-1:0] count  // count output
);

always_ff @ (posedge clk)
    if (rst) count <= {WIDTH{1'b0}};
    else if (en) count <= count + {{WIDTH-1{1'b0}}, en};
    else count <= count - {{WIDTH-1{1'b0}},1'b1};

endmodule

